
`include "dynamic_node_top_wrap.v"




module mesh (
    input clk,
    input reset_in,

    input [`DATA_WIDTH-1:0] data_in_p_0_0,
    input  valid_in_p_0_0,
    input  yummy_in_p_0_0,
    output [`DATA_WIDTH-1:0] data_out_p_0_0,
    output  valid_out_p_0_0,
    output  yummy_out_p_0_0,
    output thanks_in_p_0_0,

    input [`DATA_WIDTH-1:0] data_in_p_0_1,
    input  valid_in_p_0_1,
    input  yummy_in_p_0_1,
    output [`DATA_WIDTH-1:0] data_out_p_0_1,
    output  valid_out_p_0_1,
    output  yummy_out_p_0_1,
    output thanks_in_p_0_1,

    input [`DATA_WIDTH-1:0] data_in_p_0_2,
    input  valid_in_p_0_2,
    input  yummy_in_p_0_2,
    output [`DATA_WIDTH-1:0] data_out_p_0_2,
    output  valid_out_p_0_2,
    output  yummy_out_p_0_2,
    output thanks_in_p_0_2,

    input [`DATA_WIDTH-1:0] data_in_p_0_3,
    input  valid_in_p_0_3,
    input  yummy_in_p_0_3,
    output [`DATA_WIDTH-1:0] data_out_p_0_3,
    output  valid_out_p_0_3,
    output  yummy_out_p_0_3,
    output thanks_in_p_0_3,

    input [`DATA_WIDTH-1:0] data_in_p_0_4,
    input  valid_in_p_0_4,
    input  yummy_in_p_0_4,
    output [`DATA_WIDTH-1:0] data_out_p_0_4,
    output  valid_out_p_0_4,
    output  yummy_out_p_0_4,
    output thanks_in_p_0_4,

    input [`DATA_WIDTH-1:0] data_in_p_1_0,
    input  valid_in_p_1_0,
    input  yummy_in_p_1_0,
    output [`DATA_WIDTH-1:0] data_out_p_1_0,
    output  valid_out_p_1_0,
    output  yummy_out_p_1_0,
    output thanks_in_p_1_0,

    input [`DATA_WIDTH-1:0] data_in_p_1_1,
    input  valid_in_p_1_1,
    input  yummy_in_p_1_1,
    output [`DATA_WIDTH-1:0] data_out_p_1_1,
    output  valid_out_p_1_1,
    output  yummy_out_p_1_1,
    output thanks_in_p_1_1,

    input [`DATA_WIDTH-1:0] data_in_p_1_2,
    input  valid_in_p_1_2,
    input  yummy_in_p_1_2,
    output [`DATA_WIDTH-1:0] data_out_p_1_2,
    output  valid_out_p_1_2,
    output  yummy_out_p_1_2,
    output thanks_in_p_1_2,

    input [`DATA_WIDTH-1:0] data_in_p_1_3,
    input  valid_in_p_1_3,
    input  yummy_in_p_1_3,
    output [`DATA_WIDTH-1:0] data_out_p_1_3,
    output  valid_out_p_1_3,
    output  yummy_out_p_1_3,
    output thanks_in_p_1_3,

    input [`DATA_WIDTH-1:0] data_in_p_1_4,
    input  valid_in_p_1_4,
    input  yummy_in_p_1_4,
    output [`DATA_WIDTH-1:0] data_out_p_1_4,
    output  valid_out_p_1_4,
    output  yummy_out_p_1_4,
    output thanks_in_p_1_4,

    input [`DATA_WIDTH-1:0] data_in_p_2_0,
    input  valid_in_p_2_0,
    input  yummy_in_p_2_0,
    output [`DATA_WIDTH-1:0] data_out_p_2_0,
    output  valid_out_p_2_0,
    output  yummy_out_p_2_0,
    output thanks_in_p_2_0,

    input [`DATA_WIDTH-1:0] data_in_p_2_1,
    input  valid_in_p_2_1,
    input  yummy_in_p_2_1,
    output [`DATA_WIDTH-1:0] data_out_p_2_1,
    output  valid_out_p_2_1,
    output  yummy_out_p_2_1,
    output thanks_in_p_2_1,

    input [`DATA_WIDTH-1:0] data_in_p_2_2,
    input  valid_in_p_2_2,
    input  yummy_in_p_2_2,
    output [`DATA_WIDTH-1:0] data_out_p_2_2,
    output  valid_out_p_2_2,
    output  yummy_out_p_2_2,
    output thanks_in_p_2_2,

    input [`DATA_WIDTH-1:0] data_in_p_2_3,
    input  valid_in_p_2_3,
    input  yummy_in_p_2_3,
    output [`DATA_WIDTH-1:0] data_out_p_2_3,
    output  valid_out_p_2_3,
    output  yummy_out_p_2_3,
    output thanks_in_p_2_3,

    input [`DATA_WIDTH-1:0] data_in_p_2_4,
    input  valid_in_p_2_4,
    input  yummy_in_p_2_4,
    output [`DATA_WIDTH-1:0] data_out_p_2_4,
    output  valid_out_p_2_4,
    output  yummy_out_p_2_4,
    output thanks_in_p_2_4,

    input [`DATA_WIDTH-1:0] data_in_p_3_0,
    input  valid_in_p_3_0,
    input  yummy_in_p_3_0,
    output [`DATA_WIDTH-1:0] data_out_p_3_0,
    output  valid_out_p_3_0,
    output  yummy_out_p_3_0,
    output thanks_in_p_3_0,

    input [`DATA_WIDTH-1:0] data_in_p_3_1,
    input  valid_in_p_3_1,
    input  yummy_in_p_3_1,
    output [`DATA_WIDTH-1:0] data_out_p_3_1,
    output  valid_out_p_3_1,
    output  yummy_out_p_3_1,
    output thanks_in_p_3_1,

    input [`DATA_WIDTH-1:0] data_in_p_3_2,
    input  valid_in_p_3_2,
    input  yummy_in_p_3_2,
    output [`DATA_WIDTH-1:0] data_out_p_3_2,
    output  valid_out_p_3_2,
    output  yummy_out_p_3_2,
    output thanks_in_p_3_2,

    input [`DATA_WIDTH-1:0] data_in_p_3_3,
    input  valid_in_p_3_3,
    input  yummy_in_p_3_3,
    output [`DATA_WIDTH-1:0] data_out_p_3_3,
    output  valid_out_p_3_3,
    output  yummy_out_p_3_3,
    output thanks_in_p_3_3,

    input [`DATA_WIDTH-1:0] data_in_p_3_4,
    input  valid_in_p_3_4,
    input  yummy_in_p_3_4,
    output [`DATA_WIDTH-1:0] data_out_p_3_4,
    output  valid_out_p_3_4,
    output  yummy_out_p_3_4,
    output thanks_in_p_3_4,

    input [`DATA_WIDTH-1:0] data_in_p_4_0,
    input  valid_in_p_4_0,
    input  yummy_in_p_4_0,
    output [`DATA_WIDTH-1:0] data_out_p_4_0,
    output  valid_out_p_4_0,
    output  yummy_out_p_4_0,
    output thanks_in_p_4_0,

    input [`DATA_WIDTH-1:0] data_in_p_4_1,
    input  valid_in_p_4_1,
    input  yummy_in_p_4_1,
    output [`DATA_WIDTH-1:0] data_out_p_4_1,
    output  valid_out_p_4_1,
    output  yummy_out_p_4_1,
    output thanks_in_p_4_1,

    input [`DATA_WIDTH-1:0] data_in_p_4_2,
    input  valid_in_p_4_2,
    input  yummy_in_p_4_2,
    output [`DATA_WIDTH-1:0] data_out_p_4_2,
    output  valid_out_p_4_2,
    output  yummy_out_p_4_2,
    output thanks_in_p_4_2,

    input [`DATA_WIDTH-1:0] data_in_p_4_3,
    input  valid_in_p_4_3,
    input  yummy_in_p_4_3,
    output [`DATA_WIDTH-1:0] data_out_p_4_3,
    output  valid_out_p_4_3,
    output  yummy_out_p_4_3,
    output thanks_in_p_4_3,

    input [`DATA_WIDTH-1:0] data_in_p_4_4,
    input  valid_in_p_4_4,
    input  yummy_in_p_4_4,
    output [`DATA_WIDTH-1:0] data_out_p_4_4,
    output  valid_out_p_4_4,
    output  yummy_out_p_4_4,
    output thanks_in_p_4_4


);

    wire [`DATA_WIDTH-1:0] data_out_n_0_0;
    wire [`DATA_WIDTH-1:0] data_out_e_0_0;
    wire [`DATA_WIDTH-1:0] data_out_s_0_0;
    wire [`DATA_WIDTH-1:0] data_out_w_0_0;

    wire valid_out_n_0_0;
    wire valid_out_e_0_0;
    wire valid_out_s_0_0;
    wire valid_out_w_0_0;

    wire yummy_out_n_0_0;
    wire yummy_out_e_0_0;
    wire yummy_out_s_0_0;
    wire yummy_out_w_0_0;

    wire [`DATA_WIDTH-1:0] data_out_n_0_1;
    wire [`DATA_WIDTH-1:0] data_out_e_0_1;
    wire [`DATA_WIDTH-1:0] data_out_s_0_1;
    wire [`DATA_WIDTH-1:0] data_out_w_0_1;

    wire valid_out_n_0_1;
    wire valid_out_e_0_1;
    wire valid_out_s_0_1;
    wire valid_out_w_0_1;

    wire yummy_out_n_0_1;
    wire yummy_out_e_0_1;
    wire yummy_out_s_0_1;
    wire yummy_out_w_0_1;

    wire [`DATA_WIDTH-1:0] data_out_n_0_2;
    wire [`DATA_WIDTH-1:0] data_out_e_0_2;
    wire [`DATA_WIDTH-1:0] data_out_s_0_2;
    wire [`DATA_WIDTH-1:0] data_out_w_0_2;

    wire valid_out_n_0_2;
    wire valid_out_e_0_2;
    wire valid_out_s_0_2;
    wire valid_out_w_0_2;

    wire yummy_out_n_0_2;
    wire yummy_out_e_0_2;
    wire yummy_out_s_0_2;
    wire yummy_out_w_0_2;

    wire [`DATA_WIDTH-1:0] data_out_n_0_3;
    wire [`DATA_WIDTH-1:0] data_out_e_0_3;
    wire [`DATA_WIDTH-1:0] data_out_s_0_3;
    wire [`DATA_WIDTH-1:0] data_out_w_0_3;

    wire valid_out_n_0_3;
    wire valid_out_e_0_3;
    wire valid_out_s_0_3;
    wire valid_out_w_0_3;

    wire yummy_out_n_0_3;
    wire yummy_out_e_0_3;
    wire yummy_out_s_0_3;
    wire yummy_out_w_0_3;

    wire [`DATA_WIDTH-1:0] data_out_n_0_4;
    wire [`DATA_WIDTH-1:0] data_out_e_0_4;
    wire [`DATA_WIDTH-1:0] data_out_s_0_4;
    wire [`DATA_WIDTH-1:0] data_out_w_0_4;

    wire valid_out_n_0_4;
    wire valid_out_e_0_4;
    wire valid_out_s_0_4;
    wire valid_out_w_0_4;

    wire yummy_out_n_0_4;
    wire yummy_out_e_0_4;
    wire yummy_out_s_0_4;
    wire yummy_out_w_0_4;

    wire [`DATA_WIDTH-1:0] data_out_n_1_0;
    wire [`DATA_WIDTH-1:0] data_out_e_1_0;
    wire [`DATA_WIDTH-1:0] data_out_s_1_0;
    wire [`DATA_WIDTH-1:0] data_out_w_1_0;

    wire valid_out_n_1_0;
    wire valid_out_e_1_0;
    wire valid_out_s_1_0;
    wire valid_out_w_1_0;

    wire yummy_out_n_1_0;
    wire yummy_out_e_1_0;
    wire yummy_out_s_1_0;
    wire yummy_out_w_1_0;

    wire [`DATA_WIDTH-1:0] data_out_n_1_1;
    wire [`DATA_WIDTH-1:0] data_out_e_1_1;
    wire [`DATA_WIDTH-1:0] data_out_s_1_1;
    wire [`DATA_WIDTH-1:0] data_out_w_1_1;

    wire valid_out_n_1_1;
    wire valid_out_e_1_1;
    wire valid_out_s_1_1;
    wire valid_out_w_1_1;

    wire yummy_out_n_1_1;
    wire yummy_out_e_1_1;
    wire yummy_out_s_1_1;
    wire yummy_out_w_1_1;

    wire [`DATA_WIDTH-1:0] data_out_n_1_2;
    wire [`DATA_WIDTH-1:0] data_out_e_1_2;
    wire [`DATA_WIDTH-1:0] data_out_s_1_2;
    wire [`DATA_WIDTH-1:0] data_out_w_1_2;

    wire valid_out_n_1_2;
    wire valid_out_e_1_2;
    wire valid_out_s_1_2;
    wire valid_out_w_1_2;

    wire yummy_out_n_1_2;
    wire yummy_out_e_1_2;
    wire yummy_out_s_1_2;
    wire yummy_out_w_1_2;

    wire [`DATA_WIDTH-1:0] data_out_n_1_3;
    wire [`DATA_WIDTH-1:0] data_out_e_1_3;
    wire [`DATA_WIDTH-1:0] data_out_s_1_3;
    wire [`DATA_WIDTH-1:0] data_out_w_1_3;

    wire valid_out_n_1_3;
    wire valid_out_e_1_3;
    wire valid_out_s_1_3;
    wire valid_out_w_1_3;

    wire yummy_out_n_1_3;
    wire yummy_out_e_1_3;
    wire yummy_out_s_1_3;
    wire yummy_out_w_1_3;

    wire [`DATA_WIDTH-1:0] data_out_n_1_4;
    wire [`DATA_WIDTH-1:0] data_out_e_1_4;
    wire [`DATA_WIDTH-1:0] data_out_s_1_4;
    wire [`DATA_WIDTH-1:0] data_out_w_1_4;

    wire valid_out_n_1_4;
    wire valid_out_e_1_4;
    wire valid_out_s_1_4;
    wire valid_out_w_1_4;

    wire yummy_out_n_1_4;
    wire yummy_out_e_1_4;
    wire yummy_out_s_1_4;
    wire yummy_out_w_1_4;

    wire [`DATA_WIDTH-1:0] data_out_n_2_0;
    wire [`DATA_WIDTH-1:0] data_out_e_2_0;
    wire [`DATA_WIDTH-1:0] data_out_s_2_0;
    wire [`DATA_WIDTH-1:0] data_out_w_2_0;

    wire valid_out_n_2_0;
    wire valid_out_e_2_0;
    wire valid_out_s_2_0;
    wire valid_out_w_2_0;

    wire yummy_out_n_2_0;
    wire yummy_out_e_2_0;
    wire yummy_out_s_2_0;
    wire yummy_out_w_2_0;

    wire [`DATA_WIDTH-1:0] data_out_n_2_1;
    wire [`DATA_WIDTH-1:0] data_out_e_2_1;
    wire [`DATA_WIDTH-1:0] data_out_s_2_1;
    wire [`DATA_WIDTH-1:0] data_out_w_2_1;

    wire valid_out_n_2_1;
    wire valid_out_e_2_1;
    wire valid_out_s_2_1;
    wire valid_out_w_2_1;

    wire yummy_out_n_2_1;
    wire yummy_out_e_2_1;
    wire yummy_out_s_2_1;
    wire yummy_out_w_2_1;

    wire [`DATA_WIDTH-1:0] data_out_n_2_2;
    wire [`DATA_WIDTH-1:0] data_out_e_2_2;
    wire [`DATA_WIDTH-1:0] data_out_s_2_2;
    wire [`DATA_WIDTH-1:0] data_out_w_2_2;

    wire valid_out_n_2_2;
    wire valid_out_e_2_2;
    wire valid_out_s_2_2;
    wire valid_out_w_2_2;

    wire yummy_out_n_2_2;
    wire yummy_out_e_2_2;
    wire yummy_out_s_2_2;
    wire yummy_out_w_2_2;

    wire [`DATA_WIDTH-1:0] data_out_n_2_3;
    wire [`DATA_WIDTH-1:0] data_out_e_2_3;
    wire [`DATA_WIDTH-1:0] data_out_s_2_3;
    wire [`DATA_WIDTH-1:0] data_out_w_2_3;

    wire valid_out_n_2_3;
    wire valid_out_e_2_3;
    wire valid_out_s_2_3;
    wire valid_out_w_2_3;

    wire yummy_out_n_2_3;
    wire yummy_out_e_2_3;
    wire yummy_out_s_2_3;
    wire yummy_out_w_2_3;

    wire [`DATA_WIDTH-1:0] data_out_n_2_4;
    wire [`DATA_WIDTH-1:0] data_out_e_2_4;
    wire [`DATA_WIDTH-1:0] data_out_s_2_4;
    wire [`DATA_WIDTH-1:0] data_out_w_2_4;

    wire valid_out_n_2_4;
    wire valid_out_e_2_4;
    wire valid_out_s_2_4;
    wire valid_out_w_2_4;

    wire yummy_out_n_2_4;
    wire yummy_out_e_2_4;
    wire yummy_out_s_2_4;
    wire yummy_out_w_2_4;

    wire [`DATA_WIDTH-1:0] data_out_n_3_0;
    wire [`DATA_WIDTH-1:0] data_out_e_3_0;
    wire [`DATA_WIDTH-1:0] data_out_s_3_0;
    wire [`DATA_WIDTH-1:0] data_out_w_3_0;

    wire valid_out_n_3_0;
    wire valid_out_e_3_0;
    wire valid_out_s_3_0;
    wire valid_out_w_3_0;

    wire yummy_out_n_3_0;
    wire yummy_out_e_3_0;
    wire yummy_out_s_3_0;
    wire yummy_out_w_3_0;

    wire [`DATA_WIDTH-1:0] data_out_n_3_1;
    wire [`DATA_WIDTH-1:0] data_out_e_3_1;
    wire [`DATA_WIDTH-1:0] data_out_s_3_1;
    wire [`DATA_WIDTH-1:0] data_out_w_3_1;

    wire valid_out_n_3_1;
    wire valid_out_e_3_1;
    wire valid_out_s_3_1;
    wire valid_out_w_3_1;

    wire yummy_out_n_3_1;
    wire yummy_out_e_3_1;
    wire yummy_out_s_3_1;
    wire yummy_out_w_3_1;

    wire [`DATA_WIDTH-1:0] data_out_n_3_2;
    wire [`DATA_WIDTH-1:0] data_out_e_3_2;
    wire [`DATA_WIDTH-1:0] data_out_s_3_2;
    wire [`DATA_WIDTH-1:0] data_out_w_3_2;

    wire valid_out_n_3_2;
    wire valid_out_e_3_2;
    wire valid_out_s_3_2;
    wire valid_out_w_3_2;

    wire yummy_out_n_3_2;
    wire yummy_out_e_3_2;
    wire yummy_out_s_3_2;
    wire yummy_out_w_3_2;

    wire [`DATA_WIDTH-1:0] data_out_n_3_3;
    wire [`DATA_WIDTH-1:0] data_out_e_3_3;
    wire [`DATA_WIDTH-1:0] data_out_s_3_3;
    wire [`DATA_WIDTH-1:0] data_out_w_3_3;

    wire valid_out_n_3_3;
    wire valid_out_e_3_3;
    wire valid_out_s_3_3;
    wire valid_out_w_3_3;

    wire yummy_out_n_3_3;
    wire yummy_out_e_3_3;
    wire yummy_out_s_3_3;
    wire yummy_out_w_3_3;

    wire [`DATA_WIDTH-1:0] data_out_n_3_4;
    wire [`DATA_WIDTH-1:0] data_out_e_3_4;
    wire [`DATA_WIDTH-1:0] data_out_s_3_4;
    wire [`DATA_WIDTH-1:0] data_out_w_3_4;

    wire valid_out_n_3_4;
    wire valid_out_e_3_4;
    wire valid_out_s_3_4;
    wire valid_out_w_3_4;

    wire yummy_out_n_3_4;
    wire yummy_out_e_3_4;
    wire yummy_out_s_3_4;
    wire yummy_out_w_3_4;

    wire [`DATA_WIDTH-1:0] data_out_n_4_0;
    wire [`DATA_WIDTH-1:0] data_out_e_4_0;
    wire [`DATA_WIDTH-1:0] data_out_s_4_0;
    wire [`DATA_WIDTH-1:0] data_out_w_4_0;

    wire valid_out_n_4_0;
    wire valid_out_e_4_0;
    wire valid_out_s_4_0;
    wire valid_out_w_4_0;

    wire yummy_out_n_4_0;
    wire yummy_out_e_4_0;
    wire yummy_out_s_4_0;
    wire yummy_out_w_4_0;

    wire [`DATA_WIDTH-1:0] data_out_n_4_1;
    wire [`DATA_WIDTH-1:0] data_out_e_4_1;
    wire [`DATA_WIDTH-1:0] data_out_s_4_1;
    wire [`DATA_WIDTH-1:0] data_out_w_4_1;

    wire valid_out_n_4_1;
    wire valid_out_e_4_1;
    wire valid_out_s_4_1;
    wire valid_out_w_4_1;

    wire yummy_out_n_4_1;
    wire yummy_out_e_4_1;
    wire yummy_out_s_4_1;
    wire yummy_out_w_4_1;

    wire [`DATA_WIDTH-1:0] data_out_n_4_2;
    wire [`DATA_WIDTH-1:0] data_out_e_4_2;
    wire [`DATA_WIDTH-1:0] data_out_s_4_2;
    wire [`DATA_WIDTH-1:0] data_out_w_4_2;

    wire valid_out_n_4_2;
    wire valid_out_e_4_2;
    wire valid_out_s_4_2;
    wire valid_out_w_4_2;

    wire yummy_out_n_4_2;
    wire yummy_out_e_4_2;
    wire yummy_out_s_4_2;
    wire yummy_out_w_4_2;

    wire [`DATA_WIDTH-1:0] data_out_n_4_3;
    wire [`DATA_WIDTH-1:0] data_out_e_4_3;
    wire [`DATA_WIDTH-1:0] data_out_s_4_3;
    wire [`DATA_WIDTH-1:0] data_out_w_4_3;

    wire valid_out_n_4_3;
    wire valid_out_e_4_3;
    wire valid_out_s_4_3;
    wire valid_out_w_4_3;

    wire yummy_out_n_4_3;
    wire yummy_out_e_4_3;
    wire yummy_out_s_4_3;
    wire yummy_out_w_4_3;

    wire [`DATA_WIDTH-1:0] data_out_n_4_4;
    wire [`DATA_WIDTH-1:0] data_out_e_4_4;
    wire [`DATA_WIDTH-1:0] data_out_s_4_4;
    wire [`DATA_WIDTH-1:0] data_out_w_4_4;

    wire valid_out_n_4_4;
    wire valid_out_e_4_4;
    wire valid_out_s_4_4;
    wire valid_out_w_4_4;

    wire yummy_out_n_4_4;
    wire yummy_out_e_4_4;
    wire yummy_out_s_4_4;
    wire yummy_out_w_4_4;


    dynamic_node_top_wrap router_0_0(
        .clk(clk),
        .reset_in(reset_in),

        .myLocX(8'd0),
        .myLocY(8'd0),
        .myChipID(14'd0),

        .dataIn_N(`DATA_WIDTH'b0),
        .yummyIn_N(1'b0),
        .validIn_N(1'b0),
        .dataOut_N(),
        .yummyOut_N(),
        .validOut_N(),

        .dataIn_S(data_out_n_0_1),
        .yummyIn_S(yummy_out_n_0_1),
        .validIn_S(valid_out_n_0_1),
        .dataOut_S(data_out_s_0_0),
        .yummyOut_S(yummy_out_s_0_0),
        .validOut_S(valid_out_s_0_0),

        .dataIn_W(`DATA_WIDTH'b0),
        .yummyIn_W(1'b0),
        .validIn_W(1'b0),
        .dataOut_W(),
        .yummyOut_W(),
        .validOut_W(),

        .dataIn_E(data_out_w_1_0),
        .yummyIn_E(yummy_out_w_1_0),
        .validIn_E(valid_out_w_1_0),
        .dataOut_E(data_out_e_0_0),
        .yummyOut_E(yummy_out_e_0_0),
        .validOut_E(valid_out_e_0_0),

        .dataIn_P(data_in_p_0_0),
        .yummyIn_P(yummy_in_p_0_0),
        .validIn_P(valid_in_p_0_0),
        .dataOut_P(data_out_p_0_0),
        .yummyOut_P(yummy_out_p_0_0),
        .validOut_P(valid_out_p_0_0),

        .thanksIn_P(thanks_in_p_0_0)

    );

    dynamic_node_top_wrap router_0_1(
        .clk(clk),
        .reset_in(reset_in),

        .myLocX(8'd0),
        .myLocY(8'd1),
        .myChipID(14'd0),

        .dataIn_N(data_out_s_0_0),
        .yummyIn_N(yummy_out_s_0_0),
        .validIn_N(valid_out_s_0_0),
        .dataOut_N(data_out_n_0_1),
        .yummyOut_N(yummy_out_n_0_1),
        .validOut_N(valid_out_n_0_1),

        .dataIn_S(data_out_n_0_2),
        .yummyIn_S(yummy_out_n_0_2),
        .validIn_S(valid_out_n_0_2),
        .dataOut_S(data_out_s_0_1),
        .yummyOut_S(yummy_out_s_0_1),
        .validOut_S(valid_out_s_0_1),

        .dataIn_W(`DATA_WIDTH'b0),
        .yummyIn_W(1'b0),
        .validIn_W(1'b0),
        .dataOut_W(),
        .yummyOut_W(),
        .validOut_W(),

        .dataIn_E(data_out_w_1_1),
        .yummyIn_E(yummy_out_w_1_1),
        .validIn_E(valid_out_w_1_1),
        .dataOut_E(data_out_e_0_1),
        .yummyOut_E(yummy_out_e_0_1),
        .validOut_E(valid_out_e_0_1),

        .dataIn_P(data_in_p_0_1),
        .yummyIn_P(yummy_in_p_0_1),
        .validIn_P(valid_in_p_0_1),
        .dataOut_P(data_out_p_0_1),
        .yummyOut_P(yummy_out_p_0_1),
        .validOut_P(valid_out_p_0_1),

        .thanksIn_P(thanks_in_p_0_1)

    );

    dynamic_node_top_wrap router_0_2(
        .clk(clk),
        .reset_in(reset_in),

        .myLocX(8'd0),
        .myLocY(8'd2),
        .myChipID(14'd0),

        .dataIn_N(data_out_s_0_1),
        .yummyIn_N(yummy_out_s_0_1),
        .validIn_N(valid_out_s_0_1),
        .dataOut_N(data_out_n_0_2),
        .yummyOut_N(yummy_out_n_0_2),
        .validOut_N(valid_out_n_0_2),

        .dataIn_S(data_out_n_0_3),
        .yummyIn_S(yummy_out_n_0_3),
        .validIn_S(valid_out_n_0_3),
        .dataOut_S(data_out_s_0_2),
        .yummyOut_S(yummy_out_s_0_2),
        .validOut_S(valid_out_s_0_2),

        .dataIn_W(`DATA_WIDTH'b0),
        .yummyIn_W(1'b0),
        .validIn_W(1'b0),
        .dataOut_W(),
        .yummyOut_W(),
        .validOut_W(),

        .dataIn_E(data_out_w_1_2),
        .yummyIn_E(yummy_out_w_1_2),
        .validIn_E(valid_out_w_1_2),
        .dataOut_E(data_out_e_0_2),
        .yummyOut_E(yummy_out_e_0_2),
        .validOut_E(valid_out_e_0_2),

        .dataIn_P(data_in_p_0_2),
        .yummyIn_P(yummy_in_p_0_2),
        .validIn_P(valid_in_p_0_2),
        .dataOut_P(data_out_p_0_2),
        .yummyOut_P(yummy_out_p_0_2),
        .validOut_P(valid_out_p_0_2),

        .thanksIn_P(thanks_in_p_0_2)

    );

    dynamic_node_top_wrap router_0_3(
        .clk(clk),
        .reset_in(reset_in),

        .myLocX(8'd0),
        .myLocY(8'd3),
        .myChipID(14'd0),

        .dataIn_N(data_out_s_0_2),
        .yummyIn_N(yummy_out_s_0_2),
        .validIn_N(valid_out_s_0_2),
        .dataOut_N(data_out_n_0_3),
        .yummyOut_N(yummy_out_n_0_3),
        .validOut_N(valid_out_n_0_3),

        .dataIn_S(data_out_n_0_4),
        .yummyIn_S(yummy_out_n_0_4),
        .validIn_S(valid_out_n_0_4),
        .dataOut_S(data_out_s_0_3),
        .yummyOut_S(yummy_out_s_0_3),
        .validOut_S(valid_out_s_0_3),

        .dataIn_W(`DATA_WIDTH'b0),
        .yummyIn_W(1'b0),
        .validIn_W(1'b0),
        .dataOut_W(),
        .yummyOut_W(),
        .validOut_W(),

        .dataIn_E(data_out_w_1_3),
        .yummyIn_E(yummy_out_w_1_3),
        .validIn_E(valid_out_w_1_3),
        .dataOut_E(data_out_e_0_3),
        .yummyOut_E(yummy_out_e_0_3),
        .validOut_E(valid_out_e_0_3),

        .dataIn_P(data_in_p_0_3),
        .yummyIn_P(yummy_in_p_0_3),
        .validIn_P(valid_in_p_0_3),
        .dataOut_P(data_out_p_0_3),
        .yummyOut_P(yummy_out_p_0_3),
        .validOut_P(valid_out_p_0_3),

        .thanksIn_P(thanks_in_p_0_3)

    );

    dynamic_node_top_wrap router_0_4(
        .clk(clk),
        .reset_in(reset_in),

        .myLocX(8'd0),
        .myLocY(8'd4),
        .myChipID(14'd0),

        .dataIn_N(data_out_s_0_3),
        .yummyIn_N(yummy_out_s_0_3),
        .validIn_N(valid_out_s_0_3),
        .dataOut_N(data_out_n_0_4),
        .yummyOut_N(yummy_out_n_0_4),
        .validOut_N(valid_out_n_0_4),

        .dataIn_S(`DATA_WIDTH'b0),
        .yummyIn_S(1'b0),
        .validIn_S(1'b0),
        .dataOut_S(),
        .yummyOut_S(),
        .validOut_S(),

        .dataIn_W(`DATA_WIDTH'b0),
        .yummyIn_W(1'b0),
        .validIn_W(1'b0),
        .dataOut_W(),
        .yummyOut_W(),
        .validOut_W(),

        .dataIn_E(data_out_w_1_4),
        .yummyIn_E(yummy_out_w_1_4),
        .validIn_E(valid_out_w_1_4),
        .dataOut_E(data_out_e_0_4),
        .yummyOut_E(yummy_out_e_0_4),
        .validOut_E(valid_out_e_0_4),

        .dataIn_P(data_in_p_0_4),
        .yummyIn_P(yummy_in_p_0_4),
        .validIn_P(valid_in_p_0_4),
        .dataOut_P(data_out_p_0_4),
        .yummyOut_P(yummy_out_p_0_4),
        .validOut_P(valid_out_p_0_4),

        .thanksIn_P(thanks_in_p_0_4)

    );

    dynamic_node_top_wrap router_1_0(
        .clk(clk),
        .reset_in(reset_in),

        .myLocX(8'd1),
        .myLocY(8'd0),
        .myChipID(14'd0),

        .dataIn_N(`DATA_WIDTH'b0),
        .yummyIn_N(1'b0),
        .validIn_N(1'b0),
        .dataOut_N(),
        .yummyOut_N(),
        .validOut_N(),

        .dataIn_S(data_out_n_1_1),
        .yummyIn_S(yummy_out_n_1_1),
        .validIn_S(valid_out_n_1_1),
        .dataOut_S(data_out_s_1_0),
        .yummyOut_S(yummy_out_s_1_0),
        .validOut_S(valid_out_s_1_0),

        .dataIn_W(data_out_e_0_0),
        .yummyIn_W(yummy_out_e_0_0),
        .validIn_W(valid_out_e_0_0),
        .dataOut_W(data_out_w_1_0),
        .yummyOut_W(yummy_out_w_1_0),
        .validOut_W(valid_out_w_1_0),

        .dataIn_E(data_out_w_2_0),
        .yummyIn_E(yummy_out_w_2_0),
        .validIn_E(valid_out_w_2_0),
        .dataOut_E(data_out_e_1_0),
        .yummyOut_E(yummy_out_e_1_0),
        .validOut_E(valid_out_e_1_0),

        .dataIn_P(data_in_p_1_0),
        .yummyIn_P(yummy_in_p_1_0),
        .validIn_P(valid_in_p_1_0),
        .dataOut_P(data_out_p_1_0),
        .yummyOut_P(yummy_out_p_1_0),
        .validOut_P(valid_out_p_1_0),

        .thanksIn_P(thanks_in_p_1_0)

    );

    dynamic_node_top_wrap router_1_1(
        .clk(clk),
        .reset_in(reset_in),

        .myLocX(8'd1),
        .myLocY(8'd1),
        .myChipID(14'd0),

        .dataIn_N(data_out_s_1_0),
        .yummyIn_N(yummy_out_s_1_0),
        .validIn_N(valid_out_s_1_0),
        .dataOut_N(data_out_n_1_1),
        .yummyOut_N(yummy_out_n_1_1),
        .validOut_N(valid_out_n_1_1),

        .dataIn_S(data_out_n_1_2),
        .yummyIn_S(yummy_out_n_1_2),
        .validIn_S(valid_out_n_1_2),
        .dataOut_S(data_out_s_1_1),
        .yummyOut_S(yummy_out_s_1_1),
        .validOut_S(valid_out_s_1_1),

        .dataIn_W(data_out_e_0_1),
        .yummyIn_W(yummy_out_e_0_1),
        .validIn_W(valid_out_e_0_1),
        .dataOut_W(data_out_w_1_1),
        .yummyOut_W(yummy_out_w_1_1),
        .validOut_W(valid_out_w_1_1),

        .dataIn_E(data_out_w_2_1),
        .yummyIn_E(yummy_out_w_2_1),
        .validIn_E(valid_out_w_2_1),
        .dataOut_E(data_out_e_1_1),
        .yummyOut_E(yummy_out_e_1_1),
        .validOut_E(valid_out_e_1_1),

        .dataIn_P(data_in_p_1_1),
        .yummyIn_P(yummy_in_p_1_1),
        .validIn_P(valid_in_p_1_1),
        .dataOut_P(data_out_p_1_1),
        .yummyOut_P(yummy_out_p_1_1),
        .validOut_P(valid_out_p_1_1),

        .thanksIn_P(thanks_in_p_1_1)

    );

    dynamic_node_top_wrap router_1_2(
        .clk(clk),
        .reset_in(reset_in),

        .myLocX(8'd1),
        .myLocY(8'd2),
        .myChipID(14'd0),

        .dataIn_N(data_out_s_1_1),
        .yummyIn_N(yummy_out_s_1_1),
        .validIn_N(valid_out_s_1_1),
        .dataOut_N(data_out_n_1_2),
        .yummyOut_N(yummy_out_n_1_2),
        .validOut_N(valid_out_n_1_2),

        .dataIn_S(data_out_n_1_3),
        .yummyIn_S(yummy_out_n_1_3),
        .validIn_S(valid_out_n_1_3),
        .dataOut_S(data_out_s_1_2),
        .yummyOut_S(yummy_out_s_1_2),
        .validOut_S(valid_out_s_1_2),

        .dataIn_W(data_out_e_0_2),
        .yummyIn_W(yummy_out_e_0_2),
        .validIn_W(valid_out_e_0_2),
        .dataOut_W(data_out_w_1_2),
        .yummyOut_W(yummy_out_w_1_2),
        .validOut_W(valid_out_w_1_2),

        .dataIn_E(data_out_w_2_2),
        .yummyIn_E(yummy_out_w_2_2),
        .validIn_E(valid_out_w_2_2),
        .dataOut_E(data_out_e_1_2),
        .yummyOut_E(yummy_out_e_1_2),
        .validOut_E(valid_out_e_1_2),

        .dataIn_P(data_in_p_1_2),
        .yummyIn_P(yummy_in_p_1_2),
        .validIn_P(valid_in_p_1_2),
        .dataOut_P(data_out_p_1_2),
        .yummyOut_P(yummy_out_p_1_2),
        .validOut_P(valid_out_p_1_2),

        .thanksIn_P(thanks_in_p_1_2)

    );

    dynamic_node_top_wrap router_1_3(
        .clk(clk),
        .reset_in(reset_in),

        .myLocX(8'd1),
        .myLocY(8'd3),
        .myChipID(14'd0),

        .dataIn_N(data_out_s_1_2),
        .yummyIn_N(yummy_out_s_1_2),
        .validIn_N(valid_out_s_1_2),
        .dataOut_N(data_out_n_1_3),
        .yummyOut_N(yummy_out_n_1_3),
        .validOut_N(valid_out_n_1_3),

        .dataIn_S(data_out_n_1_4),
        .yummyIn_S(yummy_out_n_1_4),
        .validIn_S(valid_out_n_1_4),
        .dataOut_S(data_out_s_1_3),
        .yummyOut_S(yummy_out_s_1_3),
        .validOut_S(valid_out_s_1_3),

        .dataIn_W(data_out_e_0_3),
        .yummyIn_W(yummy_out_e_0_3),
        .validIn_W(valid_out_e_0_3),
        .dataOut_W(data_out_w_1_3),
        .yummyOut_W(yummy_out_w_1_3),
        .validOut_W(valid_out_w_1_3),

        .dataIn_E(data_out_w_2_3),
        .yummyIn_E(yummy_out_w_2_3),
        .validIn_E(valid_out_w_2_3),
        .dataOut_E(data_out_e_1_3),
        .yummyOut_E(yummy_out_e_1_3),
        .validOut_E(valid_out_e_1_3),

        .dataIn_P(data_in_p_1_3),
        .yummyIn_P(yummy_in_p_1_3),
        .validIn_P(valid_in_p_1_3),
        .dataOut_P(data_out_p_1_3),
        .yummyOut_P(yummy_out_p_1_3),
        .validOut_P(valid_out_p_1_3),

        .thanksIn_P(thanks_in_p_1_3)

    );

    dynamic_node_top_wrap router_1_4(
        .clk(clk),
        .reset_in(reset_in),

        .myLocX(8'd1),
        .myLocY(8'd4),
        .myChipID(14'd0),

        .dataIn_N(data_out_s_1_3),
        .yummyIn_N(yummy_out_s_1_3),
        .validIn_N(valid_out_s_1_3),
        .dataOut_N(data_out_n_1_4),
        .yummyOut_N(yummy_out_n_1_4),
        .validOut_N(valid_out_n_1_4),

        .dataIn_S(`DATA_WIDTH'b0),
        .yummyIn_S(1'b0),
        .validIn_S(1'b0),
        .dataOut_S(),
        .yummyOut_S(),
        .validOut_S(),

        .dataIn_W(data_out_e_0_4),
        .yummyIn_W(yummy_out_e_0_4),
        .validIn_W(valid_out_e_0_4),
        .dataOut_W(data_out_w_1_4),
        .yummyOut_W(yummy_out_w_1_4),
        .validOut_W(valid_out_w_1_4),

        .dataIn_E(data_out_w_2_4),
        .yummyIn_E(yummy_out_w_2_4),
        .validIn_E(valid_out_w_2_4),
        .dataOut_E(data_out_e_1_4),
        .yummyOut_E(yummy_out_e_1_4),
        .validOut_E(valid_out_e_1_4),

        .dataIn_P(data_in_p_1_4),
        .yummyIn_P(yummy_in_p_1_4),
        .validIn_P(valid_in_p_1_4),
        .dataOut_P(data_out_p_1_4),
        .yummyOut_P(yummy_out_p_1_4),
        .validOut_P(valid_out_p_1_4),

        .thanksIn_P(thanks_in_p_1_4)

    );

    dynamic_node_top_wrap router_2_0(
        .clk(clk),
        .reset_in(reset_in),

        .myLocX(8'd2),
        .myLocY(8'd0),
        .myChipID(14'd0),

        .dataIn_N(`DATA_WIDTH'b0),
        .yummyIn_N(1'b0),
        .validIn_N(1'b0),
        .dataOut_N(),
        .yummyOut_N(),
        .validOut_N(),

        .dataIn_S(data_out_n_2_1),
        .yummyIn_S(yummy_out_n_2_1),
        .validIn_S(valid_out_n_2_1),
        .dataOut_S(data_out_s_2_0),
        .yummyOut_S(yummy_out_s_2_0),
        .validOut_S(valid_out_s_2_0),

        .dataIn_W(data_out_e_1_0),
        .yummyIn_W(yummy_out_e_1_0),
        .validIn_W(valid_out_e_1_0),
        .dataOut_W(data_out_w_2_0),
        .yummyOut_W(yummy_out_w_2_0),
        .validOut_W(valid_out_w_2_0),

        .dataIn_E(data_out_w_3_0),
        .yummyIn_E(yummy_out_w_3_0),
        .validIn_E(valid_out_w_3_0),
        .dataOut_E(data_out_e_2_0),
        .yummyOut_E(yummy_out_e_2_0),
        .validOut_E(valid_out_e_2_0),

        .dataIn_P(data_in_p_2_0),
        .yummyIn_P(yummy_in_p_2_0),
        .validIn_P(valid_in_p_2_0),
        .dataOut_P(data_out_p_2_0),
        .yummyOut_P(yummy_out_p_2_0),
        .validOut_P(valid_out_p_2_0),

        .thanksIn_P(thanks_in_p_2_0)

    );

    dynamic_node_top_wrap router_2_1(
        .clk(clk),
        .reset_in(reset_in),

        .myLocX(8'd2),
        .myLocY(8'd1),
        .myChipID(14'd0),

        .dataIn_N(data_out_s_2_0),
        .yummyIn_N(yummy_out_s_2_0),
        .validIn_N(valid_out_s_2_0),
        .dataOut_N(data_out_n_2_1),
        .yummyOut_N(yummy_out_n_2_1),
        .validOut_N(valid_out_n_2_1),

        .dataIn_S(data_out_n_2_2),
        .yummyIn_S(yummy_out_n_2_2),
        .validIn_S(valid_out_n_2_2),
        .dataOut_S(data_out_s_2_1),
        .yummyOut_S(yummy_out_s_2_1),
        .validOut_S(valid_out_s_2_1),

        .dataIn_W(data_out_e_1_1),
        .yummyIn_W(yummy_out_e_1_1),
        .validIn_W(valid_out_e_1_1),
        .dataOut_W(data_out_w_2_1),
        .yummyOut_W(yummy_out_w_2_1),
        .validOut_W(valid_out_w_2_1),

        .dataIn_E(data_out_w_3_1),
        .yummyIn_E(yummy_out_w_3_1),
        .validIn_E(valid_out_w_3_1),
        .dataOut_E(data_out_e_2_1),
        .yummyOut_E(yummy_out_e_2_1),
        .validOut_E(valid_out_e_2_1),

        .dataIn_P(data_in_p_2_1),
        .yummyIn_P(yummy_in_p_2_1),
        .validIn_P(valid_in_p_2_1),
        .dataOut_P(data_out_p_2_1),
        .yummyOut_P(yummy_out_p_2_1),
        .validOut_P(valid_out_p_2_1),

        .thanksIn_P(thanks_in_p_2_1)

    );

    dynamic_node_top_wrap router_2_2(
        .clk(clk),
        .reset_in(reset_in),

        .myLocX(8'd2),
        .myLocY(8'd2),
        .myChipID(14'd0),

        .dataIn_N(data_out_s_2_1),
        .yummyIn_N(yummy_out_s_2_1),
        .validIn_N(valid_out_s_2_1),
        .dataOut_N(data_out_n_2_2),
        .yummyOut_N(yummy_out_n_2_2),
        .validOut_N(valid_out_n_2_2),

        .dataIn_S(data_out_n_2_3),
        .yummyIn_S(yummy_out_n_2_3),
        .validIn_S(valid_out_n_2_3),
        .dataOut_S(data_out_s_2_2),
        .yummyOut_S(yummy_out_s_2_2),
        .validOut_S(valid_out_s_2_2),

        .dataIn_W(data_out_e_1_2),
        .yummyIn_W(yummy_out_e_1_2),
        .validIn_W(valid_out_e_1_2),
        .dataOut_W(data_out_w_2_2),
        .yummyOut_W(yummy_out_w_2_2),
        .validOut_W(valid_out_w_2_2),

        .dataIn_E(data_out_w_3_2),
        .yummyIn_E(yummy_out_w_3_2),
        .validIn_E(valid_out_w_3_2),
        .dataOut_E(data_out_e_2_2),
        .yummyOut_E(yummy_out_e_2_2),
        .validOut_E(valid_out_e_2_2),

        .dataIn_P(data_in_p_2_2),
        .yummyIn_P(yummy_in_p_2_2),
        .validIn_P(valid_in_p_2_2),
        .dataOut_P(data_out_p_2_2),
        .yummyOut_P(yummy_out_p_2_2),
        .validOut_P(valid_out_p_2_2),

        .thanksIn_P(thanks_in_p_2_2)

    );

    dynamic_node_top_wrap router_2_3(
        .clk(clk),
        .reset_in(reset_in),

        .myLocX(8'd2),
        .myLocY(8'd3),
        .myChipID(14'd0),

        .dataIn_N(data_out_s_2_2),
        .yummyIn_N(yummy_out_s_2_2),
        .validIn_N(valid_out_s_2_2),
        .dataOut_N(data_out_n_2_3),
        .yummyOut_N(yummy_out_n_2_3),
        .validOut_N(valid_out_n_2_3),

        .dataIn_S(data_out_n_2_4),
        .yummyIn_S(yummy_out_n_2_4),
        .validIn_S(valid_out_n_2_4),
        .dataOut_S(data_out_s_2_3),
        .yummyOut_S(yummy_out_s_2_3),
        .validOut_S(valid_out_s_2_3),

        .dataIn_W(data_out_e_1_3),
        .yummyIn_W(yummy_out_e_1_3),
        .validIn_W(valid_out_e_1_3),
        .dataOut_W(data_out_w_2_3),
        .yummyOut_W(yummy_out_w_2_3),
        .validOut_W(valid_out_w_2_3),

        .dataIn_E(data_out_w_3_3),
        .yummyIn_E(yummy_out_w_3_3),
        .validIn_E(valid_out_w_3_3),
        .dataOut_E(data_out_e_2_3),
        .yummyOut_E(yummy_out_e_2_3),
        .validOut_E(valid_out_e_2_3),

        .dataIn_P(data_in_p_2_3),
        .yummyIn_P(yummy_in_p_2_3),
        .validIn_P(valid_in_p_2_3),
        .dataOut_P(data_out_p_2_3),
        .yummyOut_P(yummy_out_p_2_3),
        .validOut_P(valid_out_p_2_3),

        .thanksIn_P(thanks_in_p_2_3)

    );

    dynamic_node_top_wrap router_2_4(
        .clk(clk),
        .reset_in(reset_in),

        .myLocX(8'd2),
        .myLocY(8'd4),
        .myChipID(14'd0),

        .dataIn_N(data_out_s_2_3),
        .yummyIn_N(yummy_out_s_2_3),
        .validIn_N(valid_out_s_2_3),
        .dataOut_N(data_out_n_2_4),
        .yummyOut_N(yummy_out_n_2_4),
        .validOut_N(valid_out_n_2_4),

        .dataIn_S(`DATA_WIDTH'b0),
        .yummyIn_S(1'b0),
        .validIn_S(1'b0),
        .dataOut_S(),
        .yummyOut_S(),
        .validOut_S(),

        .dataIn_W(data_out_e_1_4),
        .yummyIn_W(yummy_out_e_1_4),
        .validIn_W(valid_out_e_1_4),
        .dataOut_W(data_out_w_2_4),
        .yummyOut_W(yummy_out_w_2_4),
        .validOut_W(valid_out_w_2_4),

        .dataIn_E(data_out_w_3_4),
        .yummyIn_E(yummy_out_w_3_4),
        .validIn_E(valid_out_w_3_4),
        .dataOut_E(data_out_e_2_4),
        .yummyOut_E(yummy_out_e_2_4),
        .validOut_E(valid_out_e_2_4),

        .dataIn_P(data_in_p_2_4),
        .yummyIn_P(yummy_in_p_2_4),
        .validIn_P(valid_in_p_2_4),
        .dataOut_P(data_out_p_2_4),
        .yummyOut_P(yummy_out_p_2_4),
        .validOut_P(valid_out_p_2_4),

        .thanksIn_P(thanks_in_p_2_4)

    );

    dynamic_node_top_wrap router_3_0(
        .clk(clk),
        .reset_in(reset_in),

        .myLocX(8'd3),
        .myLocY(8'd0),
        .myChipID(14'd0),

        .dataIn_N(`DATA_WIDTH'b0),
        .yummyIn_N(1'b0),
        .validIn_N(1'b0),
        .dataOut_N(),
        .yummyOut_N(),
        .validOut_N(),

        .dataIn_S(data_out_n_3_1),
        .yummyIn_S(yummy_out_n_3_1),
        .validIn_S(valid_out_n_3_1),
        .dataOut_S(data_out_s_3_0),
        .yummyOut_S(yummy_out_s_3_0),
        .validOut_S(valid_out_s_3_0),

        .dataIn_W(data_out_e_2_0),
        .yummyIn_W(yummy_out_e_2_0),
        .validIn_W(valid_out_e_2_0),
        .dataOut_W(data_out_w_3_0),
        .yummyOut_W(yummy_out_w_3_0),
        .validOut_W(valid_out_w_3_0),

        .dataIn_E(data_out_w_4_0),
        .yummyIn_E(yummy_out_w_4_0),
        .validIn_E(valid_out_w_4_0),
        .dataOut_E(data_out_e_3_0),
        .yummyOut_E(yummy_out_e_3_0),
        .validOut_E(valid_out_e_3_0),

        .dataIn_P(data_in_p_3_0),
        .yummyIn_P(yummy_in_p_3_0),
        .validIn_P(valid_in_p_3_0),
        .dataOut_P(data_out_p_3_0),
        .yummyOut_P(yummy_out_p_3_0),
        .validOut_P(valid_out_p_3_0),

        .thanksIn_P(thanks_in_p_3_0)

    );

    dynamic_node_top_wrap router_3_1(
        .clk(clk),
        .reset_in(reset_in),

        .myLocX(8'd3),
        .myLocY(8'd1),
        .myChipID(14'd0),

        .dataIn_N(data_out_s_3_0),
        .yummyIn_N(yummy_out_s_3_0),
        .validIn_N(valid_out_s_3_0),
        .dataOut_N(data_out_n_3_1),
        .yummyOut_N(yummy_out_n_3_1),
        .validOut_N(valid_out_n_3_1),

        .dataIn_S(data_out_n_3_2),
        .yummyIn_S(yummy_out_n_3_2),
        .validIn_S(valid_out_n_3_2),
        .dataOut_S(data_out_s_3_1),
        .yummyOut_S(yummy_out_s_3_1),
        .validOut_S(valid_out_s_3_1),

        .dataIn_W(data_out_e_2_1),
        .yummyIn_W(yummy_out_e_2_1),
        .validIn_W(valid_out_e_2_1),
        .dataOut_W(data_out_w_3_1),
        .yummyOut_W(yummy_out_w_3_1),
        .validOut_W(valid_out_w_3_1),

        .dataIn_E(data_out_w_4_1),
        .yummyIn_E(yummy_out_w_4_1),
        .validIn_E(valid_out_w_4_1),
        .dataOut_E(data_out_e_3_1),
        .yummyOut_E(yummy_out_e_3_1),
        .validOut_E(valid_out_e_3_1),

        .dataIn_P(data_in_p_3_1),
        .yummyIn_P(yummy_in_p_3_1),
        .validIn_P(valid_in_p_3_1),
        .dataOut_P(data_out_p_3_1),
        .yummyOut_P(yummy_out_p_3_1),
        .validOut_P(valid_out_p_3_1),

        .thanksIn_P(thanks_in_p_3_1)

    );

    dynamic_node_top_wrap router_3_2(
        .clk(clk),
        .reset_in(reset_in),

        .myLocX(8'd3),
        .myLocY(8'd2),
        .myChipID(14'd0),

        .dataIn_N(data_out_s_3_1),
        .yummyIn_N(yummy_out_s_3_1),
        .validIn_N(valid_out_s_3_1),
        .dataOut_N(data_out_n_3_2),
        .yummyOut_N(yummy_out_n_3_2),
        .validOut_N(valid_out_n_3_2),

        .dataIn_S(data_out_n_3_3),
        .yummyIn_S(yummy_out_n_3_3),
        .validIn_S(valid_out_n_3_3),
        .dataOut_S(data_out_s_3_2),
        .yummyOut_S(yummy_out_s_3_2),
        .validOut_S(valid_out_s_3_2),

        .dataIn_W(data_out_e_2_2),
        .yummyIn_W(yummy_out_e_2_2),
        .validIn_W(valid_out_e_2_2),
        .dataOut_W(data_out_w_3_2),
        .yummyOut_W(yummy_out_w_3_2),
        .validOut_W(valid_out_w_3_2),

        .dataIn_E(data_out_w_4_2),
        .yummyIn_E(yummy_out_w_4_2),
        .validIn_E(valid_out_w_4_2),
        .dataOut_E(data_out_e_3_2),
        .yummyOut_E(yummy_out_e_3_2),
        .validOut_E(valid_out_e_3_2),

        .dataIn_P(data_in_p_3_2),
        .yummyIn_P(yummy_in_p_3_2),
        .validIn_P(valid_in_p_3_2),
        .dataOut_P(data_out_p_3_2),
        .yummyOut_P(yummy_out_p_3_2),
        .validOut_P(valid_out_p_3_2),

        .thanksIn_P(thanks_in_p_3_2)

    );

    dynamic_node_top_wrap router_3_3(
        .clk(clk),
        .reset_in(reset_in),

        .myLocX(8'd3),
        .myLocY(8'd3),
        .myChipID(14'd0),

        .dataIn_N(data_out_s_3_2),
        .yummyIn_N(yummy_out_s_3_2),
        .validIn_N(valid_out_s_3_2),
        .dataOut_N(data_out_n_3_3),
        .yummyOut_N(yummy_out_n_3_3),
        .validOut_N(valid_out_n_3_3),

        .dataIn_S(data_out_n_3_4),
        .yummyIn_S(yummy_out_n_3_4),
        .validIn_S(valid_out_n_3_4),
        .dataOut_S(data_out_s_3_3),
        .yummyOut_S(yummy_out_s_3_3),
        .validOut_S(valid_out_s_3_3),

        .dataIn_W(data_out_e_2_3),
        .yummyIn_W(yummy_out_e_2_3),
        .validIn_W(valid_out_e_2_3),
        .dataOut_W(data_out_w_3_3),
        .yummyOut_W(yummy_out_w_3_3),
        .validOut_W(valid_out_w_3_3),

        .dataIn_E(data_out_w_4_3),
        .yummyIn_E(yummy_out_w_4_3),
        .validIn_E(valid_out_w_4_3),
        .dataOut_E(data_out_e_3_3),
        .yummyOut_E(yummy_out_e_3_3),
        .validOut_E(valid_out_e_3_3),

        .dataIn_P(data_in_p_3_3),
        .yummyIn_P(yummy_in_p_3_3),
        .validIn_P(valid_in_p_3_3),
        .dataOut_P(data_out_p_3_3),
        .yummyOut_P(yummy_out_p_3_3),
        .validOut_P(valid_out_p_3_3),

        .thanksIn_P(thanks_in_p_3_3)

    );

    dynamic_node_top_wrap router_3_4(
        .clk(clk),
        .reset_in(reset_in),

        .myLocX(8'd3),
        .myLocY(8'd4),
        .myChipID(14'd0),

        .dataIn_N(data_out_s_3_3),
        .yummyIn_N(yummy_out_s_3_3),
        .validIn_N(valid_out_s_3_3),
        .dataOut_N(data_out_n_3_4),
        .yummyOut_N(yummy_out_n_3_4),
        .validOut_N(valid_out_n_3_4),

        .dataIn_S(`DATA_WIDTH'b0),
        .yummyIn_S(1'b0),
        .validIn_S(1'b0),
        .dataOut_S(),
        .yummyOut_S(),
        .validOut_S(),

        .dataIn_W(data_out_e_2_4),
        .yummyIn_W(yummy_out_e_2_4),
        .validIn_W(valid_out_e_2_4),
        .dataOut_W(data_out_w_3_4),
        .yummyOut_W(yummy_out_w_3_4),
        .validOut_W(valid_out_w_3_4),

        .dataIn_E(data_out_w_4_4),
        .yummyIn_E(yummy_out_w_4_4),
        .validIn_E(valid_out_w_4_4),
        .dataOut_E(data_out_e_3_4),
        .yummyOut_E(yummy_out_e_3_4),
        .validOut_E(valid_out_e_3_4),

        .dataIn_P(data_in_p_3_4),
        .yummyIn_P(yummy_in_p_3_4),
        .validIn_P(valid_in_p_3_4),
        .dataOut_P(data_out_p_3_4),
        .yummyOut_P(yummy_out_p_3_4),
        .validOut_P(valid_out_p_3_4),

        .thanksIn_P(thanks_in_p_3_4)

    );

    dynamic_node_top_wrap router_4_0(
        .clk(clk),
        .reset_in(reset_in),

        .myLocX(8'd4),
        .myLocY(8'd0),
        .myChipID(14'd0),

        .dataIn_N(`DATA_WIDTH'b0),
        .yummyIn_N(1'b0),
        .validIn_N(1'b0),
        .dataOut_N(),
        .yummyOut_N(),
        .validOut_N(),

        .dataIn_S(data_out_n_4_1),
        .yummyIn_S(yummy_out_n_4_1),
        .validIn_S(valid_out_n_4_1),
        .dataOut_S(data_out_s_4_0),
        .yummyOut_S(yummy_out_s_4_0),
        .validOut_S(valid_out_s_4_0),

        .dataIn_W(data_out_e_3_0),
        .yummyIn_W(yummy_out_e_3_0),
        .validIn_W(valid_out_e_3_0),
        .dataOut_W(data_out_w_4_0),
        .yummyOut_W(yummy_out_w_4_0),
        .validOut_W(valid_out_w_4_0),

        .dataIn_E(`DATA_WIDTH'b0),
        .yummyIn_E(1'b0),
        .validIn_E(1'b0),
        .dataOut_E(),
        .yummyOut_E(),
        .validOut_E(),

        .dataIn_P(data_in_p_4_0),
        .yummyIn_P(yummy_in_p_4_0),
        .validIn_P(valid_in_p_4_0),
        .dataOut_P(data_out_p_4_0),
        .yummyOut_P(yummy_out_p_4_0),
        .validOut_P(valid_out_p_4_0),

        .thanksIn_P(thanks_in_p_4_0)

    );

    dynamic_node_top_wrap router_4_1(
        .clk(clk),
        .reset_in(reset_in),

        .myLocX(8'd4),
        .myLocY(8'd1),
        .myChipID(14'd0),

        .dataIn_N(data_out_s_4_0),
        .yummyIn_N(yummy_out_s_4_0),
        .validIn_N(valid_out_s_4_0),
        .dataOut_N(data_out_n_4_1),
        .yummyOut_N(yummy_out_n_4_1),
        .validOut_N(valid_out_n_4_1),

        .dataIn_S(data_out_n_4_2),
        .yummyIn_S(yummy_out_n_4_2),
        .validIn_S(valid_out_n_4_2),
        .dataOut_S(data_out_s_4_1),
        .yummyOut_S(yummy_out_s_4_1),
        .validOut_S(valid_out_s_4_1),

        .dataIn_W(data_out_e_3_1),
        .yummyIn_W(yummy_out_e_3_1),
        .validIn_W(valid_out_e_3_1),
        .dataOut_W(data_out_w_4_1),
        .yummyOut_W(yummy_out_w_4_1),
        .validOut_W(valid_out_w_4_1),

        .dataIn_E(`DATA_WIDTH'b0),
        .yummyIn_E(1'b0),
        .validIn_E(1'b0),
        .dataOut_E(),
        .yummyOut_E(),
        .validOut_E(),

        .dataIn_P(data_in_p_4_1),
        .yummyIn_P(yummy_in_p_4_1),
        .validIn_P(valid_in_p_4_1),
        .dataOut_P(data_out_p_4_1),
        .yummyOut_P(yummy_out_p_4_1),
        .validOut_P(valid_out_p_4_1),

        .thanksIn_P(thanks_in_p_4_1)

    );

    dynamic_node_top_wrap router_4_2(
        .clk(clk),
        .reset_in(reset_in),

        .myLocX(8'd4),
        .myLocY(8'd2),
        .myChipID(14'd0),

        .dataIn_N(data_out_s_4_1),
        .yummyIn_N(yummy_out_s_4_1),
        .validIn_N(valid_out_s_4_1),
        .dataOut_N(data_out_n_4_2),
        .yummyOut_N(yummy_out_n_4_2),
        .validOut_N(valid_out_n_4_2),

        .dataIn_S(data_out_n_4_3),
        .yummyIn_S(yummy_out_n_4_3),
        .validIn_S(valid_out_n_4_3),
        .dataOut_S(data_out_s_4_2),
        .yummyOut_S(yummy_out_s_4_2),
        .validOut_S(valid_out_s_4_2),

        .dataIn_W(data_out_e_3_2),
        .yummyIn_W(yummy_out_e_3_2),
        .validIn_W(valid_out_e_3_2),
        .dataOut_W(data_out_w_4_2),
        .yummyOut_W(yummy_out_w_4_2),
        .validOut_W(valid_out_w_4_2),

        .dataIn_E(`DATA_WIDTH'b0),
        .yummyIn_E(1'b0),
        .validIn_E(1'b0),
        .dataOut_E(),
        .yummyOut_E(),
        .validOut_E(),

        .dataIn_P(data_in_p_4_2),
        .yummyIn_P(yummy_in_p_4_2),
        .validIn_P(valid_in_p_4_2),
        .dataOut_P(data_out_p_4_2),
        .yummyOut_P(yummy_out_p_4_2),
        .validOut_P(valid_out_p_4_2),

        .thanksIn_P(thanks_in_p_4_2)

    );

    dynamic_node_top_wrap router_4_3(
        .clk(clk),
        .reset_in(reset_in),

        .myLocX(8'd4),
        .myLocY(8'd3),
        .myChipID(14'd0),

        .dataIn_N(data_out_s_4_2),
        .yummyIn_N(yummy_out_s_4_2),
        .validIn_N(valid_out_s_4_2),
        .dataOut_N(data_out_n_4_3),
        .yummyOut_N(yummy_out_n_4_3),
        .validOut_N(valid_out_n_4_3),

        .dataIn_S(data_out_n_4_4),
        .yummyIn_S(yummy_out_n_4_4),
        .validIn_S(valid_out_n_4_4),
        .dataOut_S(data_out_s_4_3),
        .yummyOut_S(yummy_out_s_4_3),
        .validOut_S(valid_out_s_4_3),

        .dataIn_W(data_out_e_3_3),
        .yummyIn_W(yummy_out_e_3_3),
        .validIn_W(valid_out_e_3_3),
        .dataOut_W(data_out_w_4_3),
        .yummyOut_W(yummy_out_w_4_3),
        .validOut_W(valid_out_w_4_3),

        .dataIn_E(`DATA_WIDTH'b0),
        .yummyIn_E(1'b0),
        .validIn_E(1'b0),
        .dataOut_E(),
        .yummyOut_E(),
        .validOut_E(),

        .dataIn_P(data_in_p_4_3),
        .yummyIn_P(yummy_in_p_4_3),
        .validIn_P(valid_in_p_4_3),
        .dataOut_P(data_out_p_4_3),
        .yummyOut_P(yummy_out_p_4_3),
        .validOut_P(valid_out_p_4_3),

        .thanksIn_P(thanks_in_p_4_3)

    );

    dynamic_node_top_wrap router_4_4(
        .clk(clk),
        .reset_in(reset_in),

        .myLocX(8'd4),
        .myLocY(8'd4),
        .myChipID(14'd0),

        .dataIn_N(data_out_s_4_3),
        .yummyIn_N(yummy_out_s_4_3),
        .validIn_N(valid_out_s_4_3),
        .dataOut_N(data_out_n_4_4),
        .yummyOut_N(yummy_out_n_4_4),
        .validOut_N(valid_out_n_4_4),

        .dataIn_S(`DATA_WIDTH'b0),
        .yummyIn_S(1'b0),
        .validIn_S(1'b0),
        .dataOut_S(),
        .yummyOut_S(),
        .validOut_S(),

        .dataIn_W(data_out_e_3_4),
        .yummyIn_W(yummy_out_e_3_4),
        .validIn_W(valid_out_e_3_4),
        .dataOut_W(data_out_w_4_4),
        .yummyOut_W(yummy_out_w_4_4),
        .validOut_W(valid_out_w_4_4),

        .dataIn_E(`DATA_WIDTH'b0),
        .yummyIn_E(1'b0),
        .validIn_E(1'b0),
        .dataOut_E(),
        .yummyOut_E(),
        .validOut_E(),

        .dataIn_P(data_in_p_4_4),
        .yummyIn_P(yummy_in_p_4_4),
        .validIn_P(valid_in_p_4_4),
        .dataOut_P(data_out_p_4_4),
        .yummyOut_P(yummy_out_p_4_4),
        .validOut_P(valid_out_p_4_4),

        .thanksIn_P(thanks_in_p_4_4)

    );




endmodule

